/*
 * FPGA Top Level for AXKU3 Ping Responder
 * Hardware: AXKU3 (XCKU3P) + FH1223 (FMC SFP)
 */
`timescale 1ns / 1ps
`default_nettype none

module fpga_top (
    // 200MHz System Clock (Bank 84)
    input  wire       sys_clk_p,
    input  wire       sys_clk_n,
    
    input  wire       rst_n, // Active Low Reset (Key)

    // SFP / GTY Interface (Bank 226 - SFP1)
    input  wire       sfp_rx_p,
    input  wire       sfp_rx_n,
    output wire       sfp_tx_p,
    output wire       sfp_tx_n,
    
    // SFP Reference Clock (From FMC - 125MHz)
    input  wire       gt_refclk_p,
    input  wire       gt_refclk_n,

    // LEDs
    output wire [3:0] led
);

    // -------------------------------------------------------------------------
    // 1. Clocking Infrastructure
    // -------------------------------------------------------------------------
    wire clk_125m;      // User logic clock from Ethernet IP (userclk2_out)
    wire clk_200m_raw;  // Output of IBUFDS
    wire clk_200m;      // Buffered system clock (Output of BUFG)
    wire clk_50m;       // DRP Clock (Generated by MMCM)
    wire mmcm_locked_sys;
    wire rst_125m;
    
    // Buffer the 200MHz System Clock from Differential Pins
    IBUFDS sys_clk_buf (.I(sys_clk_p), .IB(sys_clk_n), .O(clk_200m_raw));

    // [FIX] Insert BUFG to allow routing from IOB to MMCM in different regions
    BUFG sys_clk_global_buf (.I(clk_200m_raw), .O(clk_200m));

    // Clocking Wizard: 200MHz -> 50MHz for DRP
    // Input is now the global buffered clock (clk_200m)
    clk_wiz_0 sys_pll_inst (
        .clk_in1  (clk_200m),
        .clk_out1 (clk_50m),     // 50MHz for DRP
        .reset    (!rst_n),      // Active High Reset
        .locked   (mmcm_locked_sys)
    );

    // -------------------------------------------------------------------------
    // 2. Ethernet PCS/PMA IP (The PHY Layer)
    // -------------------------------------------------------------------------
    wire [7:0]  gmii_txd;
    wire        gmii_tx_en;
    wire        gmii_tx_er;
    wire [7:0]  gmii_rxd;
    wire        gmii_rx_dv;
    wire        gmii_rx_er;
    wire        status_link_up;
    wire        eth_mmcm_locked;
    wire [15:0] status_vector;

    // NOTE: MDIO disabled. Using configuration_vector.
    gig_ethernet_pcs_pma_0 eth_phy_inst (
        .gtrefclk_p           (gt_refclk_p),
        .gtrefclk_n           (gt_refclk_n),
        .independent_clock_bufg(clk_50m),
        
        .txp                  (sfp_tx_p),
        .txn                  (sfp_tx_n),
        .rxp                  (sfp_rx_p),
        .rxn                  (sfp_rx_n),
        
        .gmii_txd             (gmii_txd),
        .gmii_tx_en           (gmii_tx_en),
        .gmii_tx_er           (gmii_tx_er),
        .gmii_rxd             (gmii_rxd),
        .gmii_rx_dv           (gmii_rx_dv),
        .gmii_rx_er           (gmii_rx_er),
        .gmii_isolate         (),
        
        // Configuration Vector 
        // Bit 4: Auto-Neg Enable (1=Enable)
        // Bit 3: Isolate (0=Normal)
        // Bit 2: Power Down (0=Normal)
        // Bit 1: Loopback (0=Normal)
        // Bit 0: Unidirectional (0=Normal)
        .configuration_vector (5'b10000),
        
        // IMPORTANT: This port MUST be driven to avoid logic trimming errors
        // when MDIO is disabled but Auto-Negotiation is enabled.
        .an_restart_config    (1'b0), 
        .an_adv_config_vector (16'b0000000000100001), // Advertise 1000BASE-X Full Duplex (Bit 5=1, Bit 0=1)
//        .an_adv_config_val    (1'b0), // Not needed if we hold vector constant? (Actually usually needs a pulse, but let's try 0)
        
        .status_vector        (status_vector), 
        .reset                (!rst_n),
        .signal_detect        (1'b1),
        
        .mmcm_locked_out      (eth_mmcm_locked),
        .userclk_out          (),
        .userclk2_out         (clk_125m),
        .rxuserclk_out        (),
        .rxuserclk2_out       ()
    );
    
    assign status_link_up = status_vector[0];

    reg [3:0] rst_sync = 4'hF;
    always @(posedge clk_125m) rst_sync <= {rst_sync[2:0], !eth_mmcm_locked};
    assign rst_125m = rst_sync[3];

    // -------------------------------------------------------------------------
    // 3. Ethernet MAC (Verilog-Ethernet Library)
    // -------------------------------------------------------------------------
    wire [7:0]  rx_axis_tdata;
    wire        rx_axis_tvalid;
    wire        rx_axis_tlast;
    wire        rx_axis_tuser; 
    
    wire [7:0]  tx_axis_tdata;
    wire        tx_axis_tvalid;
    wire        tx_axis_tlast;
    wire        tx_axis_tready;

    eth_mac_1g #(
        .ENABLE_PADDING(1),
        .MIN_FRAME_LENGTH(10)
    ) mac_inst (        
        // Logic Interface Clocks & Resets
        .tx_clk(clk_125m),
        .tx_rst(rst_125m),
        .rx_clk(clk_125m),
        .rx_rst(rst_125m),
        
        // AXI Stream Interface
        .tx_axis_tdata(tx_axis_tdata),
        .tx_axis_tvalid(tx_axis_tvalid),
        .tx_axis_tlast(tx_axis_tlast),
        .tx_axis_tready(tx_axis_tready),
        .rx_axis_tdata(rx_axis_tdata),
        .rx_axis_tvalid(rx_axis_tvalid),
        .rx_axis_tlast(rx_axis_tlast),
        .rx_axis_tuser(rx_axis_tuser),
        
        // GMII Interface
        .gmii_rxd(gmii_rxd),
        .gmii_rx_dv(gmii_rx_dv),
        .gmii_rx_er(gmii_rx_er),
        .gmii_txd(gmii_txd),
        .gmii_tx_en(gmii_tx_en),
        .gmii_tx_er(gmii_tx_er),
        
        // Configuration
        .rx_clk_enable(1'b1),
        .tx_clk_enable(1'b1),
        .rx_mii_select(1'b0),
        .tx_mii_select(1'b0),
        // Explicit Configuration enables
        .cfg_rx_enable(1'b1), 
        .cfg_tx_enable(1'b1),
        .cfg_ifg(8'd12)
//        .cfg_rx_min_frame_length(32'd10) 
    );

    // -------------------------------------------------------------------------
    // 4. ARP Infrastructure
    // -------------------------------------------------------------------------
    
    // Signals for Ethernet Frame Extraction (RX)
    wire        rx_eth_hdr_valid;
    wire        rx_eth_hdr_ready;
    wire [47:0] rx_eth_dest_mac;
    wire [47:0] rx_eth_src_mac;
    wire [15:0] rx_eth_type;
    wire [7:0]  rx_eth_payload_axis_tdata;
    wire        rx_eth_payload_axis_tvalid;
    wire        rx_eth_payload_axis_tlast;
    wire        rx_eth_payload_axis_tuser;
    wire        rx_eth_payload_axis_tready;

    // Signals for Ethernet Frame Construction (TX)
    wire        tx_eth_hdr_valid;
    wire        tx_eth_hdr_ready;
    wire [47:0] tx_eth_dest_mac;
    wire [47:0] tx_eth_src_mac;
    wire [15:0] tx_eth_type;
    wire [7:0]  tx_eth_payload_axis_tdata;
    wire        tx_eth_payload_axis_tvalid;
    wire        tx_eth_payload_axis_tlast;
    wire        tx_eth_payload_axis_tuser;
    wire        tx_eth_payload_axis_tready;

    // RX Adapter: Raw AXI Stream (MAC) -> Split Header/Payload (ARP)
    eth_axis_rx #(
        .DATA_WIDTH(8)
    ) eth_axis_rx_inst (
        .clk(clk_125m),
        .rst(rst_125m),
        .s_axis_tdata(rx_axis_tdata),
        .s_axis_tvalid(rx_axis_tvalid),
        .s_axis_tlast(rx_axis_tlast),
        .s_axis_tuser(rx_axis_tuser),
        .s_axis_tkeep(1'b1), // [FIX] Connect Keep
        .s_axis_tready(), 
        .m_eth_hdr_valid(rx_eth_hdr_valid),
        .m_eth_hdr_ready(rx_eth_hdr_ready),
        .m_eth_dest_mac(rx_eth_dest_mac),
        .m_eth_src_mac(rx_eth_src_mac),
        .m_eth_type(rx_eth_type),
        .m_eth_payload_axis_tdata(rx_eth_payload_axis_tdata),
        .m_eth_payload_axis_tvalid(rx_eth_payload_axis_tvalid),
        .m_eth_payload_axis_tlast(rx_eth_payload_axis_tlast),
        .m_eth_payload_axis_tuser(rx_eth_payload_axis_tuser),
        .m_eth_payload_axis_tready(rx_eth_payload_axis_tready),
        .busy(),
        .error_header_early_termination()
    );

    // TX Adapter: Split Header/Payload (ARP) -> Raw AXI Stream
    wire [7:0] arp_tx_axis_tdata;
    wire       arp_tx_axis_tvalid;
    wire       arp_tx_axis_tlast;
    wire       arp_tx_axis_tready;

    eth_axis_tx #(
        .DATA_WIDTH(8)
    ) eth_axis_tx_inst (
        .clk(clk_125m),
        .rst(rst_125m),
        .s_eth_hdr_valid(tx_eth_hdr_valid),
        .s_eth_hdr_ready(tx_eth_hdr_ready),
        .s_eth_dest_mac(tx_eth_dest_mac),
        .s_eth_src_mac(tx_eth_src_mac),
        .s_eth_type(tx_eth_type),
        .s_eth_payload_axis_tdata(tx_eth_payload_axis_tdata),
        .s_eth_payload_axis_tvalid(tx_eth_payload_axis_tvalid),
        .s_eth_payload_axis_tlast(tx_eth_payload_axis_tlast),
        .s_eth_payload_axis_tuser(tx_eth_payload_axis_tuser),
        .s_eth_payload_axis_tkeep(1'b1), // [FIX] Connect Keep
        .s_eth_payload_axis_tready(tx_eth_payload_axis_tready),
        // Output as AXI Stream
        .m_axis_tdata(arp_tx_axis_tdata),
        .m_axis_tvalid(arp_tx_axis_tvalid),
        .m_axis_tlast(arp_tx_axis_tlast),
        .m_axis_tready(arp_tx_axis_tready),
        .busy()
    );

    // ARP Configuration
    localparam TARGET_IP  = {8'd192, 8'd168, 8'd1, 8'd128};
    localparam TARGET_MAC = 48'h02_00_00_00_00_00;

    // The ARP Core
    arp #(
        .DATA_WIDTH(8),
        .KEEP_ENABLE(0),
        .CACHE_ADDR_WIDTH(9)
    ) arp_inst (
        .clk(clk_125m),
        .rst(rst_125m),
        
        // Input from eth_axis_rx
        .s_eth_hdr_valid(rx_eth_hdr_valid),
        .s_eth_hdr_ready(rx_eth_hdr_ready),
        .s_eth_dest_mac(rx_eth_dest_mac),
        .s_eth_src_mac(rx_eth_src_mac),
        .s_eth_type(rx_eth_type),
        .s_eth_payload_axis_tdata(rx_eth_payload_axis_tdata),
        .s_eth_payload_axis_tkeep(1'b1), 
        .s_eth_payload_axis_tvalid(rx_eth_payload_axis_tvalid),
        .s_eth_payload_axis_tready(rx_eth_payload_axis_tready),
        .s_eth_payload_axis_tlast(rx_eth_payload_axis_tlast),
        .s_eth_payload_axis_tuser(rx_eth_payload_axis_tuser),
        
        // Output to eth_axis_tx
        .m_eth_hdr_valid(tx_eth_hdr_valid),
        .m_eth_hdr_ready(tx_eth_hdr_ready),
        .m_eth_dest_mac(tx_eth_dest_mac),
        .m_eth_src_mac(tx_eth_src_mac),
        .m_eth_type(tx_eth_type),
        .m_eth_payload_axis_tdata(tx_eth_payload_axis_tdata),
        .m_eth_payload_axis_tkeep(), 
        .m_eth_payload_axis_tvalid(tx_eth_payload_axis_tvalid),
        .m_eth_payload_axis_tready(tx_eth_payload_axis_tready),
        .m_eth_payload_axis_tlast(tx_eth_payload_axis_tlast),
        .m_eth_payload_axis_tuser(tx_eth_payload_axis_tuser),

        // ARP Logic
        .arp_request_valid(1'b0),
        .arp_request_ready(),
        .arp_request_ip(32'd0),
        .arp_response_valid(),
        .arp_response_ready(1'b1),
        .arp_response_error(),
        .arp_response_mac(),
        .local_mac(TARGET_MAC),
        .local_ip(TARGET_IP),
        .gateway_ip(32'd0),
        .subnet_mask(32'hFFFFFF00),
        .clear_cache(1'b0)
    );

    // -------------------------------------------------------------------------
    // 5. UDP Echo Engine & AXI Stream Arbiter
    // -------------------------------------------------------------------------
//    wire [7:0] icmp_tx_data;
//    wire       icmp_tx_valid, icmp_tx_last, icmp_tx_ready;
//    wire       ping_pulse;

//    icmp_echo_engine echo_inst (
//        .clk(clk_125m),
//        .rst(rst_125m),
//        .s_axis_tdata(rx_axis_tdata),   
//        .s_axis_tvalid(rx_axis_tvalid),
//        .s_axis_tlast(rx_axis_tlast),
//        .s_axis_tready(), 
//        .m_axis_tdata(icmp_tx_data),
//        .m_axis_tvalid(icmp_tx_valid),
//        .m_axis_tlast(icmp_tx_last),
//        .m_axis_tready(icmp_tx_ready),
//        .ping_detect(ping_pulse)
//    );

    wire [7:0] udp_tx_data;
    wire       udp_tx_valid, udp_tx_last, udp_tx_ready;
    wire       udp_pulse;
    
    udp_hardcoded_echo udp_inst (
        .clk(clk_125m),
        .rst(rst_125m),
        
        // RX Input
        .s_axis_tdata(rx_axis_tdata),    
        .s_axis_tvalid(rx_axis_tvalid),
        .s_axis_tlast(rx_axis_tlast),
        .s_axis_tready(), // Open or connected to logic if needed
        
        // TX Output
        .m_axis_tdata(udp_tx_data),
        .m_axis_tvalid(udp_tx_valid),
        .m_axis_tlast(udp_tx_last),
        .m_axis_tready(udp_tx_ready)
    );

    assign udp_pulse = udp_tx_valid;

    // AXI Stream Arbiter (Port 0 = UDP, Port 1 = ARP)
    axis_arb_mux #(
        .DATA_WIDTH(8),
        .S_COUNT(2),
        .ARB_TYPE_ROUND_ROBIN(1)
    ) arbiter_inst (
        .clk(clk_125m),
        .rst(rst_125m),
        
        // Output to MAC (Raw AXI Stream)
        .m_axis_tdata(tx_axis_tdata),
        .m_axis_tvalid(tx_axis_tvalid),
        .m_axis_tlast(tx_axis_tlast),
        .m_axis_tready(tx_axis_tready),
        
        // Inputs: Port 0 = UDP, Port 1 = ARP
        .s_axis_tdata({udp_tx_data, arp_tx_axis_tdata}),
        .s_axis_tvalid({udp_tx_valid, arp_tx_axis_tvalid}),
        .s_axis_tlast({udp_tx_last, arp_tx_axis_tlast}),
        .s_axis_tready({udp_tx_ready, arp_tx_axis_tready}),
        
        // Unused sideband signals
        .s_axis_tkeep(2'b11), // [FIX] Connect Keep
        .s_axis_tid(0),
        .s_axis_tdest(0),
        .s_axis_tuser(0),
        .m_axis_tkeep(),
        .m_axis_tid(),
        .m_axis_tdest(),
        .m_axis_tuser()
    );

    // -------------------------------------------------------------------------
    // 6. LED Logic
    // -------------------------------------------------------------------------
    reg [26:0] hb_cnt;
    always @(posedge clk_50m) hb_cnt <= hb_cnt + 1; 
    
    reg [23:0] ping_stretch_cnt;
    always @(posedge clk_125m) begin
        if (udp_pulse) ping_stretch_cnt <= {24{1'b1}};
        else if (ping_stretch_cnt > 0) ping_stretch_cnt <= ping_stretch_cnt - 1;
    end

    assign led[0] = hb_cnt[26];           // Heartbeat (Alive)
    assign led[1] = eth_mmcm_locked;      // Ethernet Clock Good
    assign led[2] = status_link_up;       // Link Up
    assign led[3] = |ping_stretch_cnt;    // Ping Activity
    
    // -------------------------------------------------------------------------
    // 7. Debugging (ILA)
    // -------------------------------------------------------------------------
    
    ila_0 my_ila (
        .clk(clk_125m), 
        
        // SLOT 0: RX Interface (What are we receiving?)
        .probe0(rx_axis_tdata),      // [7:0]
        .probe1(rx_axis_tvalid),     // [0:0]
        .probe2(rx_axis_tlast),      // [0:0] <-- Added
        
        // SLOT 1: TX Interface (What are we sending?)
        .probe3(tx_axis_tdata),      // [7:0]
        .probe4(tx_axis_tvalid),     // [0:0]
        .probe5(tx_axis_tlast),      // [0:0] <-- Added
        .probe6(tx_axis_tready),     // [0:0] 
        
        // SLOT 2: Internals & Status
        .probe7(udp_tx_valid),       // [0:0] <-- Tells us "It was ME who sent that!"
        .probe8(status_link_up),     // [0:0] <-- Cable status
        .probe9(eth_mmcm_locked)     // [0:0] <-- Clock status
    );

endmodule